module flash_top(
	input wire wb_clk_i
	
);

endmodule